//100KHz