//100KHz e 10KHz