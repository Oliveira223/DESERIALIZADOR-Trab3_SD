module queue(
    input logic clock,
    input logic reset,
    input logic 

);