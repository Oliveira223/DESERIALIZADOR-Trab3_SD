module queue_tb; 
