module top_module(
    input logic 
);