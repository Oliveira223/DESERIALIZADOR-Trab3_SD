//10KHz
